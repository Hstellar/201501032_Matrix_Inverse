`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Hena Ghonia 201501032
// Create Date:    10:13:39 10/07/2016 
// Design Name: 
// Module Name:    matrix inverse 
// Project Name: 

//This code does not work for floating point
//////////////////////////////////////////////////////////////////////////////////
module matrix_inverse(clk);

input clk;
real mat[0:4][0:9];

always@(posedge clk)
begin

		mat[0][0]=16'd1;   //matrix is intialized
		mat[0][1]=16'd2;
		mat[0][2]=16'd1;
		mat[0][3]=16'd0;
		mat[0][4]=16'd0;
		mat[0][5]=16'd1;
		mat[0][6]=16'd0;
		mat[0][7]=16'd0;
		mat[0][8]=16'd0;
		mat[0][9]=16'd0;
		
		mat[1][0]=16'd0;
	   mat[1][1]=16'd1;
      mat[1][2]=16'd2;
      mat[1][3]=16'd1;
      mat[1][4]=16'd0;
		mat[1][5]=16'd0;
		mat[1][6]=16'd1;
		mat[1][7]=16'd0;
		mat[1][8]=16'd0;
		mat[1][9]=16'd0;

		mat[2][0]=16'd0;
      mat[2][1]=16'd0;
		mat[2][2]=16'd1;
		mat[2][3]=16'd2;
		mat[2][4]=16'd1;
		mat[2][5]=16'd0;
		mat[2][6]=16'd0;
		mat[2][7]=16'd1;
		mat[2][8]=16'd0;
		mat[2][9]=16'd0;
		
		
		mat[3][0]=16'd0;
		mat[3][1]=16'd0;
		mat[3][2]=16'd0;
		mat[3][3]=16'd1;
		mat[3][4]=16'd2;
		mat[3][5]=16'd0;
		mat[3][6]=16'd0;
		mat[3][7]=16'd0;
		mat[3][8]=16'd1;
		mat[3][9]=16'd0;
		
		mat[4][0]=16'd0;
		mat[4][1]=16'd0;
		mat[4][2]=16'd0;
		mat[4][3]=16'd0;
		mat[4][4]=16'd1;
		mat[4][5]=16'd0;
		mat[4][6]=16'd0;
		mat[4][7]=16'd0;
		mat[4][8]=16'd0;
		mat[4][9]=16'd1;


		//1st pivot
		if(mat[0][0]!=0)
		begin
		mat[0][0]=mat[0][0]/mat[0][0];
		mat[0][1]=mat[0][1]/mat[0][0];
		mat[0][2]=mat[0][2]/mat[0][0];
		mat[0][3]=mat[0][3]/mat[0][0];
		mat[0][4]=mat[0][4]/mat[0][0];
		mat[0][5]=mat[0][5]/mat[0][0];
		mat[0][6]=mat[0][6]/mat[0][0];
		mat[0][7]=mat[0][7]/mat[0][0];
		mat[0][8]=mat[0][8]/mat[0][0];
		mat[0][9]=mat[0][9]/mat[0][0];
		
		mat[1][0]=mat[1][0]+(-mat[1][0]*mat[0][0]);
		mat[1][1]=mat[1][1]+(-mat[1][0]*mat[0][1]);
		mat[1][2]=mat[1][2]+(-mat[1][0]*mat[0][2]);
		mat[1][3]=mat[1][3]+(-mat[1][0]*mat[0][3]);
		mat[1][4]=mat[1][4]+(-mat[1][0]*mat[0][4]);
		mat[1][5]=mat[1][5]+(-mat[1][0]*mat[0][5]);
		mat[1][6]=mat[1][6]+(-mat[1][0]*mat[0][6]);
		mat[1][7]=mat[1][7]+(-mat[1][0]*mat[0][7]);
		mat[1][8]=mat[1][8]+(-mat[1][0]*mat[0][8]);
		mat[1][9]=mat[1][9]+(-mat[1][0]*mat[0][9]);
		
		
		
		
		mat[2][0]=mat[2][0]+(-mat[2][0]*mat[0][0]);
		mat[2][1]=mat[2][1]+(-mat[2][0]*mat[0][1]);
		mat[2][2]=mat[2][2]+(-mat[2][0]*mat[0][2]);
		mat[2][3]=mat[2][3]+(-mat[2][0]*mat[0][3]);
		mat[2][4]=mat[2][4]+(-mat[2][0]*mat[0][4]);
		mat[2][5]=mat[2][5]+(-mat[2][0]*mat[0][5]);
		mat[2][6]=mat[2][6]+(-mat[2][0]*mat[0][6]);
		mat[2][7]=mat[2][7]+(-mat[2][0]*mat[0][7]);
		mat[2][8]=mat[2][8]+(-mat[2][0]*mat[0][8]);
		mat[2][9]=mat[2][9]+(-mat[2][0]*mat[0][9]);
		
				
		
		mat[3][0]=mat[3][0]+(-mat[3][0]*mat[0][0]);
		mat[3][1]=mat[3][1]+(-mat[3][0]*mat[0][1]);
		mat[3][2]=mat[3][2]+(-mat[3][0]*mat[0][2]);
		mat[3][3]=mat[3][3]+(-mat[3][0]*mat[0][3]);
		mat[3][4]=mat[3][4]+(-mat[3][0]*mat[0][4]);
		mat[3][5]=mat[3][5]+(-mat[3][0]*mat[0][5]);
		mat[3][6]=mat[3][6]+(-mat[3][0]*mat[0][6]);
		mat[3][7]=mat[3][7]+(-mat[3][0]*mat[0][7]);
		mat[3][8]=mat[3][8]+(-mat[3][0]*mat[0][8]);
		mat[3][9]=mat[3][9]+(-mat[3][0]*mat[0][9]);

				
		
		mat[4][0]=mat[4][0]+(-mat[4][0]*mat[0][0]);
		mat[4][1]=mat[4][1]+(-mat[4][0]*mat[0][1]);
		mat[4][2]=mat[4][2]+(-mat[4][0]*mat[0][2]);
		mat[4][3]=mat[4][3]+(-mat[4][0]*mat[0][3]);
		mat[4][4]=mat[4][4]+(-mat[4][0]*mat[0][4]);
		mat[4][5]=mat[4][5]+(-mat[4][0]*mat[0][5]);
		mat[4][6]=mat[4][6]+(-mat[4][0]*mat[0][6]);
		mat[4][7]=mat[4][7]+(-mat[4][0]*mat[0][7]);
		mat[4][8]=mat[4][8]+(-mat[4][0]*mat[0][8]);
		mat[4][9]=mat[4][9]+(-mat[4][0]*mat[0][9]);

		end
		//2nd pivot
		if(mat[1][1]!=0)
		begin
		mat[1][0]=mat[1][0]/mat[1][1];
		mat[1][1]=mat[1][1]/mat[1][1];
		mat[1][2]=mat[1][2]/mat[1][1];
		mat[1][3]=mat[1][3]/mat[1][1];
		mat[1][4]=mat[1][4]/mat[1][1];
		mat[1][5]=mat[1][5]/mat[1][1];
		mat[1][6]=mat[1][6]/mat[1][1];
		mat[1][7]=mat[1][7]/mat[1][1];
		mat[1][8]=mat[1][8]/mat[1][1];
		mat[1][9]=mat[1][9]/mat[1][1];
		
		mat[2][0]=mat[2][0]+(-mat[2][1]*mat[1][0]);
		mat[2][1]=mat[2][1]+(-mat[2][1]*mat[1][1]);
		mat[2][2]=mat[2][2]+(-mat[2][1]*mat[1][2]);
		mat[2][3]=mat[2][3]+(-mat[2][1]*mat[1][3]);
		mat[2][4]=mat[2][4]+(-mat[2][1]*mat[1][4]);
		mat[2][5]=mat[2][5]+(-mat[2][1]*mat[1][5]);
		mat[2][6]=mat[2][6]+(-mat[2][1]*mat[1][6]);
		mat[2][7]=mat[2][7]+(-mat[2][1]*mat[1][7]);
		mat[2][8]=mat[2][8]+(-mat[2][1]*mat[1][8]);
		mat[2][9]=mat[2][9]+(-mat[2][1]*mat[1][9]);
		
		mat[3][0]=mat[3][0]+(-mat[3][1]*mat[1][0]);
		mat[3][1]=mat[3][1]+(-mat[3][1]*mat[1][1]);
		mat[3][2]=mat[3][2]+(-mat[3][1]*mat[1][2]);
		mat[3][3]=mat[3][3]+(-mat[3][1]*mat[1][3]);
		mat[3][4]=mat[3][4]+(-mat[3][1]*mat[1][4]);
		mat[3][5]=mat[3][5]+(-mat[3][1]*mat[1][5]);
		mat[3][6]=mat[3][6]+(-mat[3][1]*mat[1][6]);
		mat[3][7]=mat[3][7]+(-mat[3][1]*mat[1][7]);
		mat[3][8]=mat[3][8]+(-mat[3][1]*mat[1][8]);
		mat[3][9]=mat[3][9]+(-mat[3][1]*mat[1][9]);
	
		mat[4][0]=mat[4][0]+(-mat[4][1]*mat[1][0]);
		mat[4][1]=mat[4][1]+(-mat[4][1]*mat[1][1]);
		mat[4][2]=mat[4][2]+(-mat[4][1]*mat[1][2]);
		mat[4][3]=mat[4][3]+(-mat[4][1]*mat[1][3]);
		mat[4][4]=mat[4][4]+(-mat[4][1]*mat[1][4]);
		mat[4][5]=mat[4][5]+(-mat[4][1]*mat[1][5]);
		mat[4][6]=mat[4][6]+(-mat[4][1]*mat[1][6]);
		mat[4][7]=mat[4][7]+(-mat[4][1]*mat[1][7]);
		mat[4][8]=mat[4][8]+(-mat[4][1]*mat[1][8]);
		mat[4][9]=mat[4][9]+(-mat[4][1]*mat[1][9]);
		end
		//3rd pivot
		if(mat[2][2]!=0)
		begin
		mat[2][0]=mat[2][0]/mat[2][2];
		mat[2][1]=mat[2][1]/mat[2][2];
		mat[2][2]=mat[2][2]/mat[2][2];
		mat[2][3]=mat[2][3]/mat[2][2];
		mat[2][4]=mat[2][4]/mat[2][2];
		mat[2][5]=mat[2][5]/mat[2][2];
		mat[2][6]=mat[2][6]/mat[2][2];
		mat[2][7]=mat[2][7]/mat[2][2];
		mat[2][8]=mat[2][8]/mat[2][2];
		mat[2][9]=mat[2][9]/mat[2][2];
		
		mat[3][0]=mat[3][0]+(-mat[3][2]*mat[2][0]);
		mat[3][1]=mat[3][1]+(-mat[3][2]*mat[2][1]);
		mat[3][2]=mat[3][2]+(-mat[3][2]*mat[2][2]);
		mat[3][3]=mat[3][3]+(-mat[3][2]*mat[2][3]);
		mat[3][4]=mat[3][4]+(-mat[3][2]*mat[2][4]);
		mat[3][5]=mat[3][5]+(-mat[3][2]*mat[2][5]);
		mat[3][6]=mat[3][6]+(-mat[3][2]*mat[2][6]);
		mat[3][7]=mat[3][7]+(-mat[3][2]*mat[2][7]);
		mat[3][8]=mat[3][8]+(-mat[3][2]*mat[2][8]);
		mat[3][9]=mat[3][9]+(-mat[3][2]*mat[2][9]);
		
		mat[4][0]=mat[4][0]+(-mat[4][2]*mat[2][0]);
		mat[4][1]=mat[4][1]+(-mat[4][2]*mat[2][1]);
		mat[4][2]=mat[4][2]+(-mat[4][2]*mat[2][2]);
		mat[4][3]=mat[4][3]+(-mat[4][2]*mat[2][3]);
		mat[4][4]=mat[4][4]+(-mat[4][2]*mat[2][4]);
		mat[4][5]=mat[4][5]+(-mat[4][2]*mat[2][5]);
		mat[4][6]=mat[4][6]+(-mat[4][2]*mat[2][6]);
		mat[4][7]=mat[4][7]+(-mat[4][2]*mat[2][7]);
		mat[4][8]=mat[4][8]+(-mat[4][2]*mat[2][8]);
		mat[4][9]=mat[4][9]+(-mat[4][2]*mat[2][9]);
		end
		//4th pivot
		
		if(mat[3][3]!=0)
		begin
		mat[3][0]=mat[3][0]/mat[3][3];
		mat[3][1]=mat[3][1]/mat[3][3];
		mat[3][2]=mat[3][2]/mat[3][3];
		mat[3][3]=mat[3][3]/mat[3][3];
		mat[3][4]=mat[3][4]/mat[3][3];
		mat[3][5]=mat[3][5]/mat[3][3];
		mat[3][6]=mat[3][6]/mat[3][3];
		mat[3][7]=mat[3][7]/mat[3][3];
		mat[3][8]=mat[3][8]/mat[3][3];
		mat[3][9]=mat[3][9]/mat[3][3];
		
		mat[4][0]=mat[4][0]+(-mat[4][3]*mat[3][0]);
		mat[4][1]=mat[4][1]+(-mat[4][3]*mat[3][1]);
		mat[4][2]=mat[4][2]+(-mat[4][3]*mat[3][2]);
		mat[4][3]=mat[4][3]+(-mat[4][3]*mat[3][3]);
		mat[4][4]=mat[4][4]+(-mat[4][3]*mat[3][4]);
		mat[4][5]=mat[4][5]+(-mat[4][3]*mat[3][5]);
		mat[4][6]=mat[4][6]+(-mat[4][3]*mat[3][6]);
		mat[4][7]=mat[4][7]+(-mat[4][3]*mat[3][7]);
		mat[4][8]=mat[4][8]+(-mat[4][3]*mat[3][8]);
		mat[4][9]=mat[4][9]+(-mat[4][3]*mat[3][9]);
		end
		//5th pivot
		if(mat[4][4]!=0)
		begin
		mat[4][0]=mat[4][0]/mat[4][4];
		mat[4][1]=mat[4][1]/mat[4][4];
		mat[4][2]=mat[4][2]/mat[4][4];
		mat[4][3]=mat[4][3]/mat[4][4];
		mat[4][4]=mat[4][4]/mat[4][4];
		mat[4][5]=mat[4][5]/mat[4][4];
		mat[4][6]=mat[4][6]/mat[4][4];
		mat[4][7]=mat[4][7]/mat[4][4];
		mat[4][8]=mat[4][8]/mat[4][4];
		mat[4][9]=mat[4][9]/mat[4][4];
		end
		
		
		//2nd pivot uper
		mat[0][0]=mat[0][0]+(-mat[0][1]*mat[1][0]);
		mat[0][1]=mat[0][1]+(-mat[0][1]*mat[1][1]);
		mat[0][2]=mat[0][2]+(-mat[0][1]*mat[1][2]);
		mat[0][3]=mat[0][3]+(-mat[0][1]*mat[1][3]);
		mat[0][4]=mat[0][4]+(-mat[0][1]*mat[1][4]);
		mat[0][5]=mat[0][5]+(-mat[0][1]*mat[1][5]);
		mat[0][6]=mat[0][6]+(-mat[0][1]*mat[1][6]);
		mat[0][7]=mat[0][7]+(-mat[0][1]*mat[1][7]);
		mat[0][8]=mat[0][8]+(-mat[0][1]*mat[1][8]);
		mat[0][9]=mat[0][9]+(-mat[0][1]*mat[1][9]);
		
		//3nd pivot uper
		mat[1][0]=mat[1][0]+(-mat[1][2]*mat[2][0]);
		mat[1][1]=mat[1][1]+(-mat[1][2]*mat[2][1]);
		mat[1][2]=mat[1][2]+(-mat[1][2]*mat[2][2]);
		mat[1][3]=mat[1][3]+(-mat[1][2]*mat[2][3]);
		mat[1][4]=mat[1][4]+(-mat[1][2]*mat[2][4]);
		mat[1][5]=mat[1][5]+(-mat[1][2]*mat[2][5]);
		mat[1][6]=mat[1][6]+(-mat[1][2]*mat[2][6]);
		mat[1][7]=mat[1][7]+(-mat[1][2]*mat[2][7]);
		mat[1][8]=mat[1][8]+(-mat[1][2]*mat[2][8]);
		mat[1][9]=mat[1][9]+(-mat[1][2]*mat[2][9]);
		
		mat[0][0]=mat[0][0]+(-mat[0][2]*mat[2][0]);
		mat[0][1]=mat[0][1]+(-mat[0][2]*mat[2][1]);
		mat[0][2]=mat[0][2]+(-mat[0][2]*mat[2][2]);
		mat[0][3]=mat[0][3]+(-mat[0][2]*mat[2][3]);
		mat[0][4]=mat[0][4]+(-mat[0][2]*mat[2][4]);
		mat[0][5]=mat[0][5]+(-mat[0][2]*mat[2][5]);
		mat[0][6]=mat[0][6]+(-mat[0][2]*mat[2][6]);
		mat[0][7]=mat[0][7]+(-mat[0][2]*mat[2][7]);
		mat[0][8]=mat[0][8]+(-mat[0][2]*mat[2][8]);
		mat[0][9]=mat[0][9]+(-mat[0][2]*mat[2][9]);
		
		//4th pivot uper
		
		mat[0][0]=mat[0][0]+(-mat[0][3]*mat[3][0]);
		mat[0][1]=mat[0][1]+(-mat[0][3]*mat[3][1]);
		mat[0][2]=mat[0][2]+(-mat[0][3]*mat[3][2]);
		mat[0][3]=mat[0][3]+(-mat[0][3]*mat[3][3]);
		mat[0][4]=mat[0][4]+(-mat[0][3]*mat[3][4]);
		mat[0][5]=mat[0][5]+(-mat[0][3]*mat[3][5]);
		mat[0][6]=mat[0][6]+(-mat[0][3]*mat[3][6]);
		mat[0][7]=mat[0][7]+(-mat[0][3]*mat[3][7]);
		mat[0][8]=mat[0][8]+(-mat[0][3]*mat[3][8]);
		mat[0][9]=mat[0][9]+(-mat[0][3]*mat[3][9]);
		
		mat[1][0]=mat[1][0]+(-mat[1][3]*mat[3][0]);
		mat[1][1]=mat[1][1]+(-mat[1][3]*mat[3][1]);
		mat[1][2]=mat[1][2]+(-mat[1][3]*mat[3][2]);
		mat[1][3]=mat[1][3]+(-mat[1][3]*mat[3][3]);
		mat[1][4]=mat[1][4]+(-mat[1][3]*mat[3][4]);
		mat[1][5]=mat[1][5]+(-mat[1][3]*mat[3][5]);
		mat[1][6]=mat[1][6]+(-mat[1][3]*mat[3][6]);
		mat[1][7]=mat[1][7]+(-mat[1][3]*mat[3][7]);
		mat[1][8]=mat[1][8]+(-mat[1][3]*mat[3][8]);
		mat[1][9]=mat[1][9]+(-mat[1][3]*mat[3][9]);
		
		mat[2][0]=mat[2][0]+(-mat[2][3]*mat[3][0]);
		mat[2][1]=mat[2][1]+(-mat[2][3]*mat[3][1]);
		mat[2][2]=mat[2][2]+(-mat[2][3]*mat[3][2]);
		mat[2][3]=mat[2][3]+(-mat[2][3]*mat[3][3]);
		mat[2][4]=mat[2][4]+(-mat[2][3]*mat[3][4]);
		mat[2][5]=mat[2][5]+(-mat[2][3]*mat[3][5]);
		mat[2][6]=mat[2][6]+(-mat[2][3]*mat[3][6]);
		mat[2][7]=mat[2][7]+(-mat[2][3]*mat[3][7]);
		mat[2][8]=mat[2][8]+(-mat[2][3]*mat[3][8]);
		mat[2][9]=mat[2][9]+(-mat[2][3]*mat[3][9]);
		
		
		//5th pivot upper
		
		mat[0][0]=mat[0][0]+(-mat[0][4]*mat[4][0]);
		mat[0][1]=mat[0][1]+(-mat[0][4]*mat[4][1]);
		mat[0][2]=mat[0][2]+(-mat[0][4]*mat[4][2]);
		mat[0][3]=mat[0][3]+(-mat[0][4]*mat[4][3]);
		mat[0][4]=mat[0][4]+(-mat[0][4]*mat[4][4]);
		mat[0][5]=mat[0][5]+(-mat[0][4]*mat[4][5]);
		mat[0][6]=mat[0][6]+(-mat[0][4]*mat[4][6]);
		mat[0][7]=mat[0][7]+(-mat[0][4]*mat[4][7]);
		mat[0][8]=mat[0][8]+(-mat[0][4]*mat[4][8]);
		mat[0][9]=mat[0][9]+(-mat[0][4]*mat[4][9]);
		
		mat[1][0]=mat[1][0]+(-mat[1][4]*mat[4][0]);
		mat[1][1]=mat[1][1]+(-mat[1][4]*mat[4][1]);
		mat[1][2]=mat[1][2]+(-mat[1][4]*mat[4][2]);
		mat[1][3]=mat[1][3]+(-mat[1][4]*mat[4][3]);
		mat[1][4]=mat[1][4]+(-mat[1][4]*mat[4][4]);
		mat[1][5]=mat[1][5]+(-mat[1][4]*mat[4][5]);
		mat[1][6]=mat[1][6]+(-mat[1][4]*mat[4][6]);
		mat[1][7]=mat[1][7]+(-mat[1][4]*mat[4][7]);
		mat[1][8]=mat[1][8]+(-mat[1][4]*mat[4][8]);
		mat[1][9]=mat[1][9]+(-mat[1][4]*mat[4][9]);
		
		mat[2][0]=mat[2][0]+(-mat[2][4]*mat[4][0]);
		mat[2][1]=mat[2][1]+(-mat[2][4]*mat[4][1]);
		mat[2][2]=mat[2][2]+(-mat[2][4]*mat[4][2]);
		mat[2][3]=mat[2][3]+(-mat[2][4]*mat[4][3]);
		mat[2][4]=mat[2][4]+(-mat[2][4]*mat[4][4]);
		mat[2][5]=mat[2][5]+(-mat[2][4]*mat[4][5]);
		mat[2][6]=mat[2][6]+(-mat[2][4]*mat[4][6]);
		mat[2][7]=mat[2][7]+(-mat[2][4]*mat[4][7]);
		mat[2][8]=mat[2][8]+(-mat[2][4]*mat[4][8]);
		mat[2][9]=mat[2][9]+(-mat[2][4]*mat[4][9]);
		
		mat[3][0]=mat[3][0]+(-mat[3][4]*mat[4][0]);
		mat[3][1]=mat[3][1]+(-mat[3][4]*mat[4][1]);
		mat[3][2]=mat[3][2]+(-mat[3][4]*mat[4][2]);
		mat[3][3]=mat[3][3]+(-mat[3][4]*mat[4][3]);
		mat[3][4]=mat[3][4]+(-mat[3][4]*mat[4][4]);
		mat[3][5]=mat[3][5]+(-mat[3][4]*mat[4][5]);
		mat[3][6]=mat[3][6]+(-mat[3][4]*mat[4][6]);
		mat[3][7]=mat[3][7]+(-mat[3][4]*mat[4][7]);
		mat[3][8]=mat[3][8]+(-mat[3][4]*mat[4][8]);
		mat[3][9]=mat[3][9]+(-mat[3][4]*mat[4][9]);
		

		
		$write("%f	",mat[0][5]);
		$write("%f	",mat[0][6]);
		$write("%f	",mat[0][7]);
		$write("%f	",mat[0][8]);
		$display("%f	",mat[0][9]);
		
		$write("%f	",mat[1][5]);
		$write("%f	",mat[1][6]);
		$write("%f	",mat[1][7]);
		$write("%f	",mat[1][8]);
		$display("%f	",mat[1][9]);
		
		$write("%f	",mat[2][5]);
		$write("%f	",mat[2][6]);
		$write("%f	",mat[2][7]);
		$write("%f	",mat[2][8]);
		$display("%f	",mat[2][9]);
		
		$write("%f	",mat[3][5]);
		$write("%f	",mat[3][6]);
		$write("%f	",mat[3][7]);
		$write("%f	",mat[3][8]);
		$display("%f	",mat[3][9]);
		
		$write("%f	",mat[4][5]);
		$write("%f	",mat[4][6]);
		$write("%f	",mat[4][7]);
		$write("%f	",mat[4][8]);
		$display("%f	",mat[4][9]);
		
		
		/*$write("1.0000    ");
		$write("-2.0000   ");
		$write("3.0000    ");
		$write("-4.0000   ");
		$display("5.0000		");
		
		$write("0.0000    ");
		$write("1.0000    ");
		$write("-2.0000   ");
		$write("3.0000    ");
		$display("-4.0000		");
		
		$write("0.0000    ");
		$write("0.0000    ");
		$write("1.0000    ");
		$write("-2.0000   ");
		$display("3.0000  ");

		$write("0.0000    ");
		$write("0.0000    ");
		$write("0.0000    ");
		$write("1.0000    ");
		$display("-2.0000 ");
		
		$write("0.0000    ");
		$write("0.0000    ");
		$write("0.0000    ");
		$write("0.0000    ");
		$display("1.0000");
		*/
		
end

endmodule
